`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:05:51 05/28/2015 
// Design Name: 
// Module Name:    inst_pointer_IP 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module inst_pointer_IP(
    input freeze,
    input rst,
    input clk,
    output [7:0] pc
    );


endmodule
